module q2wire(input a,b, output  y);
 
  assign y = a&b; 
endmodule
