module q4();
  reg [7:0] a = 8'b10101010;
  initial begin
    $display("a = %b",a);
  end
endmodule
