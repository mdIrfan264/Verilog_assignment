module q2reg(input a,b, output reg y);
 
  
  initial begin
    y = a&b;
 
     
     end
endmodule
