module q5();
  integer i=-5;
 
  initial begin 
    $display("i = %d",i);
    
  end
endmodule
